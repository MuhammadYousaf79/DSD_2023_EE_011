module led_circuit_comb_tb;

	logic [1:0]a1;
	logic [1:0]b1;
	logic r1;
	logic g1;
	logic be1;

led_circuit_comb uut(
.a(a1),
.b(b1),
.r(r1),
.g(g1),
.be(be1)
);

initial
begin

	a1[0] = 0; a1[1] = 0; b1[0] = 0; b1[1] = 0;
	#10;

	a1[0] = 0; a1[1] = 0; b1[0] = 0; b1[1] = 1;
	#10;

	a1[0] = 0; a1[1] = 0; b1[0] = 1; b1[1] = 0;
	#10;

	a1[0] = 0; a1[1] = 0; b1[0] = 1; b1[1] = 1;
	#10;

	a1[0] = 0; a1[1] = 1; b1[0] = 0; b1[1] = 0;
	#10;

	a1[0] = 0; a1[1] = 1; b1[0] = 0; b1[1] = 1;
	#10;

	a1[0] = 0; a1[1] = 1; b1[0] = 1; b1[1] = 0;
	#10;

	a1[0] = 0; a1[1] = 1; b1[0] = 1; b1[1] = 1;
	#10;

	a1[0] = 1; a1[1] = 0; b1[0] = 0; b1[1] = 0;
	#10;

	a1[0] = 1; a1[1] = 0; b1[0] = 0; b1[1] = 1;
	#10;

	a1[0] = 1; a1[1] = 0; b1[0] = 1; b1[1] = 0;
	#10;

	a1[0] = 1; a1[1] = 0; b1[0] = 1; b1[1] = 1;
	#10;

	a1[0] = 1; a1[1] = 1; b1[0] = 0; b1[1] = 0;
	#10;

	a1[0] = 1; a1[1] = 1; b1[0] = 0; b1[1] = 1;
	#10;

	a1[0] = 1; a1[1] = 1; b1[0] = 1; b1[1] = 0;
	#10;

	a1[0] = 1; a1[1] = 1; b1[0] = 1; b1[1] = 1;
	#10;
	$stop;
end

initial
begin
	$monitor("a0= %d, a1= %d, b0= %d, b1= %d, r= %d, g= %d, b= %d", a1[0],a1[1],b1[0],b1[1],r1,g1,be1);
end

endmodule